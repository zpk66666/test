module test
#(
parameter WIDTH = 10
)
(
input a,
output b
);
assign a = b;
endmodule